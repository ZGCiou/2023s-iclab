../00_TESTBED/TESTBED_OS.sv