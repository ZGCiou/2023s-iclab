../00_TESTBED/PATTERN_OS.sv