../00_TESTBED/TESTBED_bridge.sv