../02_SYN/Netlist/bridge_Wrapper.sv