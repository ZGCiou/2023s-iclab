../00_TESTBED/PATTERN_bridge.sv