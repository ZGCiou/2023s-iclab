../02_SYN/Netlist/OS_Wrapper.sv