../00_TESTBED/Usertype_OS.sv